`timescale 1ns / 1ps

/// \brief Template interface for VeSPA Custom Bus slave device
/// \input i_Clk Source Clock signal for the slave device, logic is processed on rising edges of this signal
/// \input i_Rst Reset signal for the device, active high
/// \input i_WEnable Write Enable signal. If this signal is set to high during a rising edge of the clock,
/// data is writen to the slave register file
/// \input i_WAddr Address of the register file that data should be writen to. This is a virtual address,
/// that should be generated by a Bus Interconnect device
/// \input i_WData Data writen to the slave register file if all the required conditions are complied
/// \input i_REnable Read Enable signal. If this signal is set to high during a rising edge of the clock,
/// data is read from the slave register file
/// \input i_RAddr Address of the register file that data will be read from. Simmilar to the i_WAddr, this
/// address should be generated by a Bus Interconnect device
/// \output o_RData When a read operation occurs, data is put on this output
/// \output o_Err This signal indicated an internal error occured on the device, such as an invalid address
module SlaveInterface
(
    //Bus related signals
    input i_Clk,
    input i_Rst,
    input i_WEnable,
    input [31:0] i_WAddr,
    input [31:0] i_WData,
    input i_REnable,
    input [31:0] i_RAddr,
    output reg [31:0] o_RData,
    output reg o_Err
    //User signals begin here
);

//Change this according to the needs of your slave
parameter REGFILE_SIZE = 4;

reg [31:0] r_SlaveRegisterFile [(REGFILE_SIZE - 1):0];

integer i;

always @(posedge i_Clk) begin
    if (i_Rst) begin
        //Zero-out the slave register file on reset
        for (i = 0; i < REGFILE_SIZE; i = i + 1) begin
            r_SlaveRegisterFile[i] <= 0;
        end
        o_Err <= 0;
    end
    else begin
        //Check if there is a write request pending
        if (i_WEnable) begin
            //Verify it the write address is within range
            if (i_WAddr < REGFILE_SIZE) begin
                //Add any extra write logic here, i.e. write protection
                r_SlaveRegisterFile[i_WAddr] = i_WData;
                o_Err <= 0;
            end
            else begin
                o_Err <= 1;
            end
        end
        //Check if there is a read request pending
        else if (i_REnable) begin
            //Verify it the read address is within range
            if (i_RAddr < REGFILE_SIZE) begin
                //Add any extra read logic here, i.e. read clamping
                o_RData = r_SlaveRegisterFile[i_RAddr];
                o_Err <= 0;
            end
            else begin
                o_Err <= 1;
            end
        end
        else begin
            r_SlaveRegisterFile[i_WAddr] <= i_WData;
            //Do nothing
        end


    end
end


endmodule
